/***********************************************************************************************/
/*********************************  MIPS 5-stage pipeline implementation ***********************/
/***********************************************************************************************/

module cpu(input clock, input reset);
 reg [31:0] PC; 
 reg [31:0] IFID_PCplus4,IDEX_PCplus4;
 reg [31:0] IFID_instr;
 reg [31:0] IDEX_rdA, IDEX_rdB, IDEX_signExtend;
 reg [4:0]  IDEX_instr_rt, IDEX_instr_rs, IDEX_instr_rd;                            
 reg        IDEX_RegDst, IDEX_ALUSrc;
 reg [1:0]  IDEX_ALUcntrl;
 reg        IDEX_Branch, IDEX_MemRead, IDEX_MemWrite; 
 reg        IDEX_MemToReg, IDEX_RegWrite;                
 reg [4:0]  EXMEM_RegWriteAddr, EXMEM_instr_rd; 
 reg [31:0] EXMEM_ALUOut;
 reg        EXMEM_Zero;
 reg [31:0] EXMEM_MemWriteData;
 reg        EXMEM_Branch, EXMEM_MemRead, EXMEM_MemWrite, EXMEM_RegWrite, EXMEM_MemToReg;
 reg [31:0] MEMWB_DMemOut;
 reg [4:0]  MEMWB_RegWriteAddr, MEMWB_instr_rd; 
 reg [31:0] MEMWB_ALUOut;
 reg        MEMWB_MemToReg, MEMWB_RegWrite;               
 wire [31:0] instr, ALUInA, ALUInB, ALUOut, rdA, rdB, signExtend, DMemOut, wRegData, PCIncr;
 wire Zero, RegDst, MemRead, MemWrite, MemToReg, ALUSrc, RegWrite, Branch;
 wire [5:0] opcode, func;
 wire [4:0] instr_rs, instr_rt, instr_rd, RegWriteAddr;
 wire [3:0] ALUOp;
 wire [1:0] ALUcntrl;
 wire [15:0] imm;

 reg [5:0] IDEX_Sa;
 wire  pc_write, ifid_write ,bubble_idex,bubble_ifid,bubble_exmem ;
 wire [1:0] bypassA,bypassB;
 wire [31:0] forwardA,forwardB ;
 wire [5:0] sa ; 
reg [5:0] IDEX_opcode, EXMEM_opcode;

wire [31:0] jump_or_pc ,pc_new ; 
wire [31:0] branch_adr;
reg [31:0] EXMEM_branch_adr ; 
wire PCSrc;
wire Jump_sign;
wire [31:0] jump ; 
wire Zero_add;

assign jump_or_pc = (Jump_sign)? jump : PC + 4;

assign pc_new = (PCSrc)? EXMEM_branch_adr : jump_or_pc ;

/***************** Instruction Fetch Unit (IF)  ****************/
 always @(posedge clock or negedge reset)
  begin 
    if (reset == 1'b0)     
       PC <= -1;     
    else if (PC == -1)
       PC <= 0;
    else if (pc_write == 1)
       PC <= pc_new;
  end
  
  // IFID pipeline register
 always @(posedge clock or negedge reset)
  begin 
    if (reset == 1'b0)     
      begin
	  
       IFID_PCplus4 <= 32'b0;    
       IFID_instr <= 32'b0;
    end 
    else if (ifid_write == 1'b1 && bubble_ifid == 0 )
      begin
       IFID_PCplus4 <= PC + 32'd4;
       IFID_instr <= instr;
    end
	else if ( bubble_ifid == 1 )
	begin
		IFID_instr <= 0; 
	end 
  end
  
// Instruction memory 1KB
Memory cpu_IMem(clock, reset, 1'b1, 1'b0, PC>>2, 32'b0, instr);
  
  
  
  
  
/***************** Instruction Decode Unit (ID)  ****************/
assign opcode = IFID_instr[31:26];
assign jump[25:0] = (IFID_instr[25:0]<<2);

assign jump[31:26] = 0; 
assign func = IFID_instr[5:0];
assign instr_rs = IFID_instr[25:21];
assign instr_rt = IFID_instr[20:16];
assign instr_rd = IFID_instr[15:11];
assign imm = IFID_instr[15:0];
assign signExtend = {{16{imm[15]}}, imm};
assign sa = IFID_instr [10:6];
// Register file
RegFile cpu_regs(clock, reset, instr_rs, instr_rt, MEMWB_RegWriteAddr, MEMWB_RegWrite, wRegData, rdA, rdB);

  // IDEX pipeline register
 always @(posedge clock or negedge reset)
  begin 
    if (reset == 1'b0)
      begin
       IDEX_rdA <= 32'b0;    
       IDEX_rdB <= 32'b0;
       IDEX_signExtend <= 32'b0;
       IDEX_instr_rd <= 5'b0;
       IDEX_instr_rs <= 5'b0;
       IDEX_instr_rt <= 5'b0;
       IDEX_RegDst <= 1'b0;
       IDEX_ALUcntrl <= 2'b0;
       IDEX_ALUSrc <= 1'b0;
       IDEX_Branch <= 1'b0;
       IDEX_MemRead <= 1'b0;
       IDEX_MemWrite <= 1'b0;
       IDEX_MemToReg <= 1'b0;                  
       IDEX_RegWrite <= 1'b0;
	   IDEX_opcode <= 6'b0;
    end 
    else if (bubble_idex == 0)
      begin
       IDEX_rdA <= rdA;
       IDEX_rdB <= rdB;
	   IDEX_PCplus4 <= IFID_PCplus4;
       IDEX_signExtend <= signExtend;
       IDEX_instr_rd <= instr_rd;
       IDEX_instr_rs <= instr_rs;
       IDEX_instr_rt <= instr_rt;
       IDEX_RegDst <= RegDst;
       IDEX_ALUcntrl <= ALUcntrl;
       IDEX_ALUSrc <= ALUSrc;
       IDEX_Branch <= Branch;
       IDEX_MemRead <= MemRead;
       IDEX_MemWrite <= MemWrite;
       IDEX_MemToReg <= MemToReg;                  
       IDEX_RegWrite <= RegWrite;
	   IDEX_Sa <= sa;
	   IDEX_opcode <= opcode;
    end 
	else if (bubble_idex == 1 )
	  begin 
       IDEX_RegDst <= 1'b0;
       IDEX_ALUcntrl <= 2'b0;
       IDEX_ALUSrc <= 1'b0;
       IDEX_MemRead <= 1'b0;
       IDEX_MemWrite <= 1'b0;
       IDEX_MemToReg <= 1'b0;                  
       IDEX_RegWrite <= 1'b0;
	   IDEX_Branch <= 1'b0;
	   
	  end 
	   
end 

// Main Control Unit 
control_main control_main (RegDst,
                  Branch,
                  MemRead,
                  MemWrite,
                  MemToReg,
                  ALUSrc,
                  RegWrite,
                  ALUcntrl,
				  Jump_sign,
                  opcode);
                  
// Instantiation of Control Unit that generates stalls goes here

stall stall( pc_write, ifid_write, PCSrc, instr_rs, instr_rt, IDEX_MemRead, IDEX_instr_rt,bubble_idex,bubble_exmem,bubble_ifid,Jump_sign);


                           
/***************** Execution Unit (EX)  ****************/
                 

  ALU add_alu(branch_adr,Zero_add,IDEX_PCplus4,IDEX_signExtend << 2,4'b0010);

//  ALU
ALU  #(32) cpu_alu(ALUOut, Zero, ALUInA, ALUInB, ALUOp);

assign RegWriteAddr = (IDEX_RegDst==1'b0) ? IDEX_instr_rt : IDEX_instr_rd;

 // EXMEM pipeline register
 always @(posedge clock or negedge reset)
  begin 
    if (reset == 1'b0 )     
      begin
       EXMEM_ALUOut <= 32'b0;    
       EXMEM_RegWriteAddr <= 5'b0;
       EXMEM_MemWriteData <= 32'b0;
       EXMEM_Zero <= 1'b0;
       EXMEM_Branch <= 1'b0;
       EXMEM_MemRead <= 1'b0;
       EXMEM_MemWrite <= 1'b0;
       EXMEM_MemToReg <= 1'b0;                  
       EXMEM_RegWrite <= 1'b0;
	   EXMEM_opcode <= 6'b0;
      end 
    else if (bubble_exmem == 0)
      begin 
	  
	   EXMEM_branch_adr <= branch_adr;
       EXMEM_ALUOut <= ALUOut;    
       EXMEM_RegWriteAddr <= RegWriteAddr;
       EXMEM_MemWriteData <= forwardB;//IDEX_rdB ;
       EXMEM_Zero <= Zero;
       EXMEM_Branch <= IDEX_Branch;
       EXMEM_MemRead <= IDEX_MemRead;
       EXMEM_MemWrite <= IDEX_MemWrite;
       EXMEM_MemToReg <= IDEX_MemToReg;                  
       EXMEM_RegWrite <= IDEX_RegWrite;
	   EXMEM_opcode <= IDEX_opcode;
      end
	  else if (bubble_exmem == 1 )
	  begin 
	    EXMEM_Zero <= 1'b0;
       EXMEM_Branch <= 1'b0;
       EXMEM_MemRead <= 1'b0;
       EXMEM_MemWrite <= 1'b0;
       EXMEM_MemToReg <= 1'b0;                  
       EXMEM_RegWrite <= 1'b0;
	   end 
  end
  
  // ALU control
  control_alu control_alu(ALUOp, IDEX_ALUcntrl, IDEX_signExtend[5:0]);
  
   // Instantiation of control logic for Forwarding goes here
  
  
  assign ALUInA = ( ALUOp == 4'b1000) ? IDEX_Sa : forwardA ;
  
  
  assign forwardA = (bypassA == 2'b10 ) ?  EXMEM_ALUOut :
				  (bypassA == 2'b01 ) ?  wRegData :
				  (bypassA == 2'b00 ) ?  IDEX_rdA :
				  'bx;
  
  assign  forwardB  = (bypassB == 2'b10 ) ?  EXMEM_ALUOut :
				     (bypassB == 2'b01 ) ?  wRegData :
				     (bypassB == 2'b00 ) ?  IDEX_rdB :
					 'bx;
					 
  
  assign ALUInB = (IDEX_ALUSrc == 1'b0) ? forwardB : IDEX_signExtend;
   
  
 
  
   control_bypass_ex  bypass_ex( bypassA, bypassB, IDEX_instr_rs, IDEX_instr_rt, EXMEM_RegWriteAddr,MEMWB_RegWriteAddr,EXMEM_RegWrite,MEMWB_RegWrite);
  
/***************** Memory Unit (MEM)  ****************/  

// Data memory 1KB
Memory cpu_DMem(clock, reset, EXMEM_MemRead, EXMEM_MemWrite, EXMEM_ALUOut, EXMEM_MemWriteData, DMemOut);

// MEMWB pipeline register
 always @(posedge clock or negedge reset)
  begin 
    if (reset == 1'b0)     
      begin
       MEMWB_DMemOut <= 32'b0;    
       MEMWB_ALUOut <= 32'b0;
       MEMWB_RegWriteAddr <= 5'b0;
       MEMWB_MemToReg <= 1'b0;                  
       MEMWB_RegWrite <= 1'b0;
      end 
    else 
      begin
       MEMWB_DMemOut <= DMemOut;
       MEMWB_ALUOut <= EXMEM_ALUOut;
       MEMWB_RegWriteAddr <= EXMEM_RegWriteAddr;
       MEMWB_MemToReg <= EXMEM_MemToReg;                  
       MEMWB_RegWrite <= EXMEM_RegWrite;
      end
  end

  
  PCsrc pssrc(clock ,reset,EXMEM_opcode,EXMEM_Zero,EXMEM_Branch,PCSrc);
  

/***************** WriteBack Unit (WB)  ****************/  
assign wRegData = (MEMWB_MemToReg == 1'b0) ? MEMWB_ALUOut : MEMWB_DMemOut;


endmodule
